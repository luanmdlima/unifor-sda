library verilog;
use verilog.vl_types.all;
entity operational_vlg_vec_tst is
end operational_vlg_vec_tst;
