-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
-- Created on Tue Dec 06 20:20:36 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY controller IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        c : IN STD_LOGIC := '0';
        tot_lt_s : IN STD_LOGIC := '0';
        d : OUT STD_LOGIC;
        tot_ld : OUT STD_LOGIC;
        tot_clr : OUT STD_LOGIC
    );
END controller;

ARCHITECTURE BEHAVIOR OF controller IS
    TYPE type_fstate IS (begining,waiting,add,provide,wait_not_c);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,c,tot_lt_s)
    BEGIN
        IF (reset='0') THEN
            reg_fstate <= begining;
            d <= '0';
            tot_ld <= '0';
            tot_clr <= '0';
        ELSE
            d <= '0';
            tot_ld <= '0';
            tot_clr <= '0';
            CASE fstate IS
                WHEN begining =>
                    reg_fstate <= waiting;

                    tot_ld <= '0';

                    d <= '0';

                    tot_clr <= '1';
                WHEN waiting =>
                    IF (((c = '0') AND (tot_lt_s = '0'))) THEN
                        reg_fstate <= provide;
                    ELSIF ((c = '1')) THEN
                        reg_fstate <= add;
                    ELSIF (((c = '0') AND (tot_lt_s = '1'))) THEN
                        reg_fstate <= waiting;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= waiting;
                    END IF;

                    tot_ld <= '0';

                    d <= '0';

                    tot_clr <= '0';
                WHEN add =>
                    reg_fstate <= wait_not_c;

                    tot_ld <= '1';

                    d <= '0';

                    tot_clr <= '0';
                WHEN provide =>
                    reg_fstate <= begining;

                    tot_ld <= '0';

                    d <= '1';

                    tot_clr <= '0';
                WHEN wait_not_c =>
                    IF ((c = '1')) THEN
                        reg_fstate <= wait_not_c;
                    ELSIF ((c = '0')) THEN
                        reg_fstate <= waiting;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= wait_not_c;
                    END IF;
                WHEN OTHERS => 
                    d <= 'X';
                    tot_ld <= 'X';
                    tot_clr <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
