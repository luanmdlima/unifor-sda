library verilog;
use verilog.vl_types.all;
entity counter_bcd_up_vlg_sample_tst is
    port(
        in_1            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end counter_bcd_up_vlg_sample_tst;
