-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
-- Created on Tue Dec 06 17:25:34 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY controller IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        counter : IN STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
        red : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        yellow : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        green : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        reset_counter : OUT STD_LOGIC
    );
END controller;

ARCHITECTURE BEHAVIOR OF controller IS
    TYPE type_fstate IS (state3,state4,state6,state5,state2,state1);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,counter)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            red <= "000";
            yellow <= "000";
            green <= "000";
            reset_counter <= '0';
        ELSE
            red <= "000";
            yellow <= "000";
            green <= "000";
            reset_counter <= '0';
            CASE fstate IS
                WHEN state3 =>
                    IF ((counter(4 DOWNTO 0) = "01100")) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    green <= "010";

                    yellow <= "000";

                    red <= "101";
                WHEN state4 =>
                    IF ((counter(4 DOWNTO 0) = "01110")) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    green <= "000";

                    yellow <= "010";

                    red <= "101";
                WHEN state6 =>
                    IF ((counter(4 DOWNTO 0) = "10101")) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;

                    green <= "000";

                    yellow <= "001";

                    red <= "110";
                WHEN state5 =>
                    IF ((counter(4 DOWNTO 0) = "10011")) THEN
                        reg_fstate <= state6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    green <= "001";

                    yellow <= "000";

                    red <= "110";
                WHEN state2 =>
                    IF ((counter(4 DOWNTO 0) = "00111")) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    green <= "000";

                    yellow <= "100";

                    red <= "011";
                WHEN state1 =>
                    IF ((counter(4 DOWNTO 0) = "00101")) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    IF ((counter(4 DOWNTO 0) = "10101")) THEN
                        reset_counter <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reset_counter <= '0';
                    END IF;

                    green <= "100";

                    yellow <= "000";

                    red <= "011";
                WHEN OTHERS => 
                    red <= "XXX";
                    yellow <= "XXX";
                    green <= "XXX";
                    reset_counter <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
