library verilog;
use verilog.vl_types.all;
entity funcoes_vlg_check_tst is
    port(
        s1              : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end funcoes_vlg_check_tst;
