library verilog;
use verilog.vl_types.all;
entity counter_5bit_vlg_vec_tst is
end counter_5bit_vlg_vec_tst;
