library verilog;
use verilog.vl_types.all;
entity counter_bin_n_vlg_vec_tst is
end counter_bin_n_vlg_vec_tst;
