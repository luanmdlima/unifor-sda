library verilog;
use verilog.vl_types.all;
entity system_vlg_check_tst is
    port(
        d               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end system_vlg_check_tst;
