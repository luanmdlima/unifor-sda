library verilog;
use verilog.vl_types.all;
entity mux16to1_vlg_vec_tst is
end mux16to1_vlg_vec_tst;
