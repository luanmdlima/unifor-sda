library verilog;
use verilog.vl_types.all;
entity counter_bcd_down_vlg_vec_tst is
end counter_bcd_down_vlg_vec_tst;
