library verilog;
use verilog.vl_types.all;
entity operational_vlg_check_tst is
    port(
        tot_lt_s        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end operational_vlg_check_tst;
