library verilog;
use verilog.vl_types.all;
entity semaphore_state_machine_vlg_vec_tst is
end semaphore_state_machine_vlg_vec_tst;
