library verilog;
use verilog.vl_types.all;
entity semaphore_vlg_vec_tst is
end semaphore_vlg_vec_tst;
