library verilog;
use verilog.vl_types.all;
entity funcoes_vlg_vec_tst is
end funcoes_vlg_vec_tst;
