library verilog;
use verilog.vl_types.all;
entity binary_up_down_counter_vlg_vec_tst is
end binary_up_down_counter_vlg_vec_tst;
