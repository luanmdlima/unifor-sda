library verilog;
use verilog.vl_types.all;
entity system_2_vlg_vec_tst is
end system_2_vlg_vec_tst;
