library verilog;
use verilog.vl_types.all;
entity adder_8b_vlg_vec_tst is
end adder_8b_vlg_vec_tst;
